package chip_env_pkg;

    import uvm_pkg::*;

    `include "chip_env.sv"

endpackage : chip_env_pkg